package shared_package;

bit test_finished ;
integer error_count ;
integer correct_count ;

endpackage